(* blackbox *)
module GATE(
  input  wire I1,
  input  wire I2,
  output wire O
);

endmodule
