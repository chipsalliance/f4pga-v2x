(* CLASS="input" *)
module IPAD(inpad);
    output wire inpad;

endmodule
