module CHILD(
    input  wire I,
    output wire O
);

endmodule
