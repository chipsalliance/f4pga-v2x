/*
 * Copyright 2020-2022 F4PGA Authors
 *
 * Licensed under the Apache License, Version 2.0 (the "License");
 * you may not use this file except in compliance with the License.
 * You may obtain a copy of the License at
 *
 *     http://www.apache.org/licenses/LICENSE-2.0
 *
 * Unless required by applicable law or agreed to in writing, software
 * distributed under the License is distributed on an "AS IS" BASIS,
 * WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
 * See the License for the specific language governing permissions and
 * limitations under the License.
 *
 * SPDX-License-Identifier: Apache-2.0
 */

`include "./not/not.sim.v"

(* MODES="PASSTHROUGH;INVERT" *)
module INV(I, O);
    input  wire I;
    output wire O;

    parameter MODE="PASSTHROUGH";

    // Passthrough (no inversion) mode
    generate if (MODE == "PASSTHROUGH") begin
        assign O = I;

    // Inversion with placeable inverter
    end else if (MODE == "INVERT") begin
        NOT inverter(I, O);

    end endgenerate
endmodule
