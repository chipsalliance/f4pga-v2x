/*
 * Copyright (C) 2020  The SymbiFlow Authors.
 *
 * Use of this source code is governed by a ISC-style
 * license that can be found in the LICENSE file or at
 * https://opensource.org/licenses/ISC
 */

`include "./child/child.sim.v"

module PARENT(
    input  wire I,
    output wire O
);

    wire hop1 = I;

    CHILD child (
    .I(hop1),
    .O(O)
    );

endmodule
