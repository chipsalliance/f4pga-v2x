/*
 * Copyright (C) 2020  The SymbiFlow Authors.
 *
 * Permission to use, copy, modify, and/or distribute this software for any
 * purpose with or without fee is hereby granted, provided that the above
 * copyright notice and this permission notice appear in all copies.
 *
 * THE SOFTWARE IS PROVIDED "AS IS" AND THE AUTHOR DISCLAIMS ALL WARRANTIES
 * WITH REGARD TO THIS SOFTWARE INCLUDING ALL IMPLIED WARRANTIES OF
 * MERCHANTABILITY AND FITNESS. IN NO EVENT SHALL THE AUTHOR BE LIABLE FOR
 * ANY SPECIAL, DIRECT, INDIRECT, OR CONSEQUENTIAL DAMAGES OR ANY DAMAGES
 * WHATSOEVER RESULTING FROM LOSS OF USE, DATA OR PROFITS, WHETHER IN AN
 * ACTION OF CONTRACT, NEGLIGENCE OR OTHER TORTIOUS ACTION, ARISING OUT OF
 * OR IN CONNECTION WITH THE USE OR PERFORMANCE OF THIS SOFTWARE.
 */

`default_nettype none
`include "cblock/cblock.sim.v"

module CARRY (
	I0,
	I1,
	O0,
	O1,
	CIN,
	COUT
);
	input wire [3:0] I0;
	input wire [3:0] I1;

	output wire O0;
	output wire O1;

	// Implicit carry pins
	input wire CIN;
	output wire COUT;

	// Carry between the two blocks
	wire c;

	CBLOCK cblock0 (.I(I0), .O(O0), .CIN(CIN), .COUT(c));
	CBLOCK cblock1 (.I(I1), .O(O1), .CIN(c), .COUT(COUT));

endmodule
