(* blackbox *)
module FF(
  (* CLOCK *)
  input  wire CLK,
  input  wire D,
  output wire Q
);

endmodule
