(* CLASS="output" *)
module OPAD(outpad);
    input  wire outpad;

endmodule
