/*
 * Copyright (C) 2020  The SymbiFlow Authors.
 *
 * Permission to use, copy, modify, and/or distribute this software for any
 * purpose with or without fee is hereby granted, provided that the above
 * copyright notice and this permission notice appear in all copies.
 *
 * THE SOFTWARE IS PROVIDED "AS IS" AND THE AUTHOR DISCLAIMS ALL WARRANTIES
 * WITH REGARD TO THIS SOFTWARE INCLUDING ALL IMPLIED WARRANTIES OF
 * MERCHANTABILITY AND FITNESS. IN NO EVENT SHALL THE AUTHOR BE LIABLE FOR
 * ANY SPECIAL, DIRECT, INDIRECT, OR CONSEQUENTIAL DAMAGES OR ANY DAMAGES
 * WHATSOEVER RESULTING FROM LOSS OF USE, DATA OR PROFITS, WHETHER IN AN
 * ACTION OF CONTRACT, NEGLIGENCE OR OTHER TORTIOUS ACTION, ARISING OUT OF
 * OR IN CONNECTION WITH THE USE OR PERFORMANCE OF THIS SOFTWARE.
 */

`default_nettype none

(* whitebox *)
module CBLOCK (
	I,
	O,
	CIN,
	COUT
);
	input wire [3:0] I;
	(* carry="C" *)
	input wire CIN;

	(* DELAY_MATRIX_I="30e-12 30e-12 30e-12 30e-12" *)
	(* DELAY_CONST_CIN="30e-12" *)
	output wire O;

	(* carry="C" *)
	(* DELAY_MATRIX_I="30e-12 30e-12 30e-12 30e-12" *)
	(* DELAY_CONST_CIN="30e-12" *)
	output wire COUT;

	wire [4:0] internal_sum;

	assign internal_sum = I + CIN;
	assign O = internal_sum[4];
	assign COUT = internal_sum[3];
endmodule
