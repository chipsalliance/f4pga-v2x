/*
 * Copyright (C) 2020  The SymbiFlow Authors.
 *
 * Use of this source code is governed by a ISC-style
 * license that can be found in the LICENSE file or at
 * https://opensource.org/licenses/ISC
 *
 * SPDX-License-Identifier:	ISC
 */

(* whitebox *)
module INPUT_NAMED_REGEX(
    input  wire clk,
    input  wire Clk,
    input  wire CLK,
    input  wire clkX,
    input  wire clkBus,
    input  wire sys_clk,
    input  wire sys_clk10,
    input  wire regular_input,
    output wire o
);

endmodule
